// Author: N/A
// Source: N/A
module maj3(input[0:2] x, f);
  maj(f, x[0], x[1], x[2]);
endmodule
